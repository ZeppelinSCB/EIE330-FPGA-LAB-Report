module SimpleVGADisplay


endmodule