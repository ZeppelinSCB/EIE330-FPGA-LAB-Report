module clk_gen(
    input wire sys_clk, // System clock, frequency is 50M Hz
    input wire sys_rst_n


    output wire locked //Check whether the phase-locked loop is locked.
);



endmodule